module memory(
    input [7:0] din,
    input [7:0] addr,
    input clk, we, 
    output [7:0] dout
);
    reg [7:0] mem_reg[15:0];
endmodule