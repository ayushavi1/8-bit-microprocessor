module memory(
    input [7:0] din,
    input [7:0] addr,
    input clk, we, 
    output [7:0] dout
);
    reg [7:0] mem_reg[255:0];

    initial
    begin
        // Assembly Code

        // Move Register Values
        mem_reg[8'h00]<=8'b0010_00_01;
        mem_reg[8'h01]<=8'b0011_10_00;
        mem_reg[8'h02]<=8'b0011_00_00;

        // Add 2 Numbers
		// mem_reg[8'h00]<=8'b0010_00_01;
		// mem_reg[8'h01]<=8'b0010_01_01;
		// mem_reg[8'h02]<=8'b0100_00_01;
		// mem_reg[8'h03]<=8'b0011_00_00;

        // Add with immediate
        // mem_reg[8'h00]<=8'b0010_00_01;
        // mem_reg[8'h01]<=8'b1100_00_01;
        // mem_reg[8'h02]<=8'b0011_00_00;

        // Subtract 2 Numbers
        // mem_reg[8'h00]<=8'b0010_00_01;
        // mem_reg[8'h01]<=8'b0010_01_11;
        // mem_reg[8'h02]<=8'b0101_00_01;
        // mem_reg[8'h03]<=8'b0011_00_00;
        
        // Subtract with immediate
        // mem_reg[8'h00]<=8'b0010_00_01;
        // mem_reg[8'h01]<=8'b1101_00_01;
        // mem_reg[8'h02]<=8'b0011_00_00;
    end

    always @(posedge clk)
	begin
		if (we)
			mem_reg[addr] <= din;
	end
	
	assign dout = mem_reg[addr];
endmodule