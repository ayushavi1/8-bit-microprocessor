module microprocessor(
    input wire ,
    output reg
);
    wire buffer;
    
endmodule