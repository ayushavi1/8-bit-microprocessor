module microcomputer(
    
);
endmodule